module up(); 

